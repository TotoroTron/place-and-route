
module top_level
#(
    parameter DATA_WIDTH = 24,
    parameter FIR_DEPTH = 128
)(
    input wire i_clk,
    input wire i_rst,
    input wire i_en,
    input wire i_din,
    input wire i_din_valid,
    output wire o_dout,
    output wire o_dout_valid
);

    wire [DATA_WIDTH-1:0] fir_din = { (LENGHT){1'b0} };
    wire [DATA_WIDTH-1:0] fir_dout = { (LENGHT){1'b0} };
    wire des_out_valid = 1'b0;
    wire fir_out_valid = 1'b0;
    wire ser_out_valid = 1'b0;

    deserializer
    #(
        .LENGTH(DATA_WIDTH)
    ) deserializer_inst (
        .i_clk(i_clk),
        .i_rst(i_rst),
        .i_en(i_en),
        .i_din(i_din),
        .i_din_valid(i_din_valid),
        .ov_dout(fir_input),
        .o_dout_valid(ser_out_valid)
    );

    fir_filter
    #(
        .DATA_WIDTH(DATA_WIDTH),
        .FIR_DEPTH(FIR_DEPTH)
    ) fir_filter_inst (
        .i_clk(i_clk),
        .i_rst(i_rst),
        .i_en(ser_out_valid),
        .iv_din(fir_din),
        .ov_dout(fir_dout),
        .o_dout_valid(fir_out_valid)
    );

    serializer
    #(
        .LENGTH(DATA_WIDTH)
    ) serializer_inst (
        .i_clk(i_clk),
        .i_rst(i_rst),
        .i_en(i_en),
        .i_din_valid(fir_out_valid),
        .i_din(fir_dout),
        .o_dout(o_dout),
        .o_dout_valid(ser_out_valid)
    );

endmodule
